library IEEE;
use IEEE.STD_LOGIC_1164.all;

ENTITY asigandorus IS
PORT(   w0, w1, w2, w3, w4 : out std_logic_vector(31 DOWNTO 0));
END asigandorus;

ARCHITECTURE synth OF asigandorus IS
BEGIN

	w0<= "00000001001000110000000100100011";
	w1<= "00010010001101000001001000110100";
	w2<= "00000001001000110100010101100111";
	w3<= "00010011000100110001001100010011";
	w4<= "00000000000000000000000000000011";


END synth;